/* CPU - top level module */

module cpu(
  input clk,
);

  always @(posedge clk) begin
    
  end

endmodule
