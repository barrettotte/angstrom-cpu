/* RAM - 12-bit addressing, 4-bit word */

module ram()



endmodule
